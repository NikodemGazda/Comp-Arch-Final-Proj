module top_tb;

// uncomment each test as needed

// `include "ram_tb.sv"
// ram_tb tb_ram();

// `include "register_tb.sv"
// register_tb tb_register();

`include "delay_tb.sv"
delay_tb tb_register();

endmodule