module top_tb;

// uncomment each test as needed

// `include "ram_tb.sv"
// ram_tb test();

// `include "register_tb.sv"
// register_tb test();

// `include "delay_tb.sv"
// delay_tb test();

`include "cache_data_tb.sv"
cache_data_tb test();

endmodule